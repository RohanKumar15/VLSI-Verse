package AHB_APB_pkg;

        import uvm_pkg::*;
        `include "uvm_macros.svh"
        `include "ahb_xtns.sv"
        `include "ahb_config.sv"
        `include "apb_config.sv"
        `include "AHB_APB_env_config.sv"
        `include "ahb_driver.sv"
        `include "ahb_monitor.sv"
        `include "ahb_sequencer.sv"
        `include "ahb_agent.sv"
        `include "ahb_agt_top.sv"
        `include "ahb_seqs.sv"

        `include "apb_xtns.sv"
        `include "apb_driver.sv"
        `include "apb_monitor.sv"
        `include "apb_sequencer.sv"
        `include "apb_agent.sv"
        `include "apb_agt_top.sv"
        `include "apb_seqs.sv"

        `include "virtual_sequencer.sv"
        `include "virtual_sequence.sv"
        `include "scoreboard.sv"

        `include "AHB_APB_env.sv"
        `include "test.sv"

endpackage
